package router_stimulus_pkg;

import uvm_pkg::*;

`include "packet.sv"
`include "packet_sequence.sv"

endpackage
